module hex

const (
	table         = '0123456789ABCDEF'
	reverse_table = [u8(0xff), 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0x00, 0x01, 0x02, 0x03, 0x04, 0x05, 0x06, 0x07, 0x08,
		0x09, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0x0a, 0x0b, 0x0c, 0x0d, 0x0e, 0x0f, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0x0a, 0x0b, 0x0c, 0x0d, 0x0e,
		0x0f, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff, 0xff,
		0xff, 0xff, 0xff, 0xff]
)

// encode_bytes converts the source bytes to hexadecimal bytes
pub fn encode_bytes(src []u8) []u8 {
	mut encoded_bytes := []u8{cap: src.len * 2}
	for val in src {
		encoded_bytes << hex.table[val >> 4]
		encoded_bytes << hex.table[val & 0x0F]
	}
	return encoded_bytes
}

// encode converts the source string into a hexadecimal string
[inline]
pub fn encode(src string) string {
	return encode_bytes(src.bytes()).bytestr()
}

// decode_bytes converts hexadecimal source bytes back into normal bytes
pub fn decode_bytes(src []u8) ![]u8 {
	if src.len % 2 != 0 {
		return error('fn hex.decode_bytes: source bytes must be divisilble by two.')
	}

	mut decoded_bytes := []u8{cap: src.len / 2}
	for i := 1; i < src.len; i += 2 {
		p := src[i - 1]
		q := src[i]

		a := hex.reverse_table[p]
		b := hex.reverse_table[q]

		if a > 0x0f {
			return error('fn hex.decode_bytes: invalid byte ${p}')
		}
		if b > 0x0f {
			return error('fn hex.decode_bytes: invalid byte ${q}')
		}
		decoded_bytes << (a << 4) | b
	}
	return decoded_bytes
}

// decode converts a hexadecimal string back into a normal string
[inline]
pub fn decode(src string) !string {
	return (decode_bytes(src.bytes())!).bytestr()
}

// encode_struct converts a struct to hexadecimal bytes
pub fn encode_struct<T>(@struct &T) ![]u8 {
	size := int(sizeof(T))
	bytes := unsafe { voidptr(@struct).vbytes(size) }
	
	if size <= 0 {
		return error('fn hex.encode_struct: struct size of zero bytes')
	}

	return encode(bytes.bytestr()).bytes()
}

// decode_struct converts hexadecimal bytes to a struct
pub fn decode_struct<T>(src []u8) !T {
	size := int(sizeof(T))
	if size <= 0 {
		return error('fn hex.decode_struct: struct size of zero bytes')
	}
	if size != src.len / 2 {
		return error('fn hex.decode_struct: struct size does not match source bytes size')
	}

	bytes := decode(src.bytestr())!
	return unsafe { *&T(bytes.bytes().data)}
}